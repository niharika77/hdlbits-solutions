//For each bit in a 32-bit vector, capture when the input signal changes from 1 in one clock cycle to 0 the next. "Capture" means
//that the output will remain 1 until the register is reset (synchronous reset).

//Each output bit behaves like a SR flip-flop: The output bit should be set (to 1) the cycle after a 1 to 0 transition 
//occurs. The output bit should be reset (to 0) at the positive clock edge when reset is high. If both of the above events 
//occur at the same time, reset has precedence. In the last 4 
//cycles of the example waveform below, the 'reset' event occurs one cycle earlier than the 'set' event, so there is no conflict here.



module top_module (
    input clk,
    input reset,
    input [31:0] in,
    output [31:0] out
);
    reg [31:0]temp;
    
    always @(posedge clk)
        begin
            temp <= in;
        end
    
    wire [31:0] temp_out;
    
    assign temp_out = temp & (~in);  // bit changing from 1 to 0
    
    reg count;
    
    always @(posedge clk)
        begin
            if(reset) begin
                count <= 0;
                out <= 0;
            end
            else 
                begin
                    if(temp_out!=0)
                    out <= temp_out;
                    else
                        out<=out;
                    end
                
        end
                        
    

endmodule
